----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:46:01 04/07/2014 
-- Design Name: 
-- Module Name:    Banco_EX - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY Banco_EX IS
	PORT (
		clk : IN STD_LOGIC;
		reset : IN STD_LOGIC;
		load : IN STD_LOGIC;
		busA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		busB : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		busA_EX : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		busB_EX : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		RegDst_ID : IN STD_LOGIC;
		ALUSrc_ID : IN STD_LOGIC;
		MemWrite_ID : IN STD_LOGIC;
		MemRead_ID : IN STD_LOGIC;
		MemtoReg_ID : IN STD_LOGIC;
		RegWrite_ID : IN STD_LOGIC;
		inm_ext : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		inm_ext_EX : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		RegDst_EX : OUT STD_LOGIC;
		ALUSrc_EX : OUT STD_LOGIC;
		MemWrite_EX : OUT STD_LOGIC;
		MemRead_EX : OUT STD_LOGIC;
		MemtoReg_EX : OUT STD_LOGIC;
		RegWrite_EX : OUT STD_LOGIC;
		-- Nuevo
		Reg_Rs_ID : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		Reg_Rs_EX : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		--Fin nuevo
		ALUctrl_ID : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		ALUctrl_EX : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		Reg_Rt_ID : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		Reg_Rd_ID : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		Reg_Rt_EX : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		Reg_Rd_EX : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		-- Nuevo excepci�n
		PC_exception_ID : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		PC_exception_EX : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		--bits de validez
		valid_I_EX_in : IN STD_LOGIC;
		valid_I_EX : OUT STD_LOGIC);
END Banco_EX;

ARCHITECTURE Behavioral OF Banco_EX IS

BEGIN
	SYNC_PROC : PROCESS (clk)
	BEGIN
		IF (clk'event AND clk = '1') THEN
			IF (reset = '1') THEN
				busA_EX <= x"00000000";
				busB_EX <= x"00000000";
				inm_ext_EX <= x"00000000";
				RegDst_EX <= '0';
				ALUSrc_EX <= '0';
				MemWrite_EX <= '0';
				MemRead_EX <= '0';
				MemtoReg_EX <= '0';
				RegWrite_EX <= '0';
				-- Nuevo
				Reg_Rs_EX <= "00000";
				PC_exception_EX <= x"00000000";
				-- fin Nuevo
				Reg_Rt_EX <= "00000";
				Reg_Rd_EX <= "00000";
				ALUctrl_EX <= "000";
				valid_I_EX <= '0';
			ELSE
				IF (load = '1') THEN
					busA_EX <= busA;
					busB_EX <= busB;
					RegDst_EX <= RegDst_ID;
					ALUSrc_EX <= ALUSrc_ID;
					MemWrite_EX <= MemWrite_ID;
					MemRead_EX <= MemRead_ID;
					MemtoReg_EX <= MemtoReg_ID;
					RegWrite_EX <= RegWrite_ID;
					-- Nuevo
					Reg_Rs_EX <= Reg_Rs_ID;
					PC_exception_EX <= PC_exception_ID;
					-- fin Nuevo
					Reg_Rt_EX <= Reg_Rt_ID;
					Reg_Rd_EX <= Reg_Rd_ID;
					ALUctrl_EX <= ALUctrl_ID;
					inm_ext_EX <= inm_ext;
					valid_I_EX <= valid_I_EX_in;
				END IF;
			END IF;
		END IF;
	END PROCESS;

END Behavioral;